module alu(
  input         reset       ,
  input         clk         ,
  input  [19:0] alu_op      ,
  input  [31:0] alu_src1    ,
  input  [31:0] alu_src2    ,
  output [31:0] alu_result  ,
  output [31:0] alu_result2 ,
  output  reg   div_ready   ,
  output  reg   result_ready,
  output        result_valid,
  output        result_valid_n
);


wire [63:0] result_data;
wire [63:0] result_data_n;
reg     dend_valid;
reg     dend_valid_n;
reg [31:0] dend_data;
reg [31:0] dend_data_n;
reg     sor_valid;
reg     sor_valid_n;
reg [31:0] sor_data;
reg [31:0] sor_data_n;
mydiv mydiv(
    .aclk           (clk            ),
    .s_axis_dividend_tvalid       (dend_valid         ),
    .s_axis_dividend_tready       (dend_ready         ),
    .s_axis_dividend_tdata        (dend_data          ),
    //被除数
    .s_axis_divisor_tvalid        (sor_valid          ),
    .s_axis_divisor_tready        (sor_ready          ),
    .s_axis_divisor_tdata         (sor_data           ),
    //除数
    .m_axis_dout_tvalid           (result_valid       ),
    .m_axis_dout_tdata            (result_data        )
);

mydiv_n mydiv_n(
    .aclk           (clk            ),
    .s_axis_dividend_tvalid       (dend_valid_n         ),
    .s_axis_dividend_tready       (dend_ready_n         ),
    .s_axis_dividend_tdata        (dend_data_n          ),
    //被除数
    .s_axis_divisor_tvalid        (sor_valid_n          ),
    .s_axis_divisor_tready        (sor_ready_n          ),
    .s_axis_divisor_tdata         (sor_data_n           ),
    //除数
    .m_axis_dout_tvalid           (result_valid_n       ),
    .m_axis_dout_tdata            (result_data_n        )
);
wire op_div;
wire op_div_n;

always @(posedge clk) begin
  if (reset) begin
    div_ready<=1;
    result_ready<=1;
  end
  if (op_div & div_ready) begin
    dend_data<=alu_src1;
    sor_data<=alu_src2;
    dend_valid<=1;
    sor_valid<=1;
    result_ready<=0;
  end
  if (op_div_n & div_ready) begin
    dend_data_n<=alu_src1;
    sor_data_n<=alu_src2;
    dend_valid_n<=1;
    sor_valid_n<=1;
    result_ready<=0;
  end
  if(dend_valid==1&dend_ready==1 &sor_valid==1&sor_ready==1) begin
    dend_valid<=0;
    sor_valid<=0;
    div_ready<=0;
    result_ready<=0;
  end
  if(dend_valid_n==1&dend_ready_n==1 &sor_valid_n==1&sor_ready_n==1) begin
    dend_valid_n<=0;
    sor_valid_n<=0;
    div_ready<=0;
    result_ready<=0;
  end
  if (result_valid_n) begin
    div_ready<=1;
    result_ready<=1;
  end
  if (result_valid) begin
    div_ready<=1;
    result_ready<=1;
  end
end


wire op_add;   //�ӷ�����
wire op_sub;   //��������
wire op_slt;   //�з��űȽϣ�С����λ
wire op_sltu;  //�޷��űȽϣ�С����λ
wire op_and;   //��λ��
wire op_nor;   //��λ���?
wire op_or;    //��λ��
wire op_xor;   //��λ���?
wire op_sll;   //�߼�����
wire op_srl;   //�߼�����
wire op_sra;   //��������
wire op_lui;   //���������ڸ߰벿��
wire op_mul;
wire op_mul_n;

assign op_add  = alu_op[ 0];
assign op_sub  = alu_op[ 1];
assign op_slt  = alu_op[ 2];
assign op_sltu = alu_op[ 3];
assign op_and  = alu_op[ 4];
assign op_nor  = alu_op[ 5];
assign op_or   = alu_op[ 6];
assign op_xor  = alu_op[ 7];
assign op_sll  = alu_op[ 8];
assign op_srl  = alu_op[ 9];
assign op_sra  = alu_op[10];
assign op_lui  = alu_op[11];
assign op_mul  = alu_op[12];
assign op_mul_n= alu_op[13];
assign op_div  = alu_op[18];
assign op_div_n= alu_op[19];

wire [31:0] add_sub_result; 
wire [31:0] slt_result; 
wire [31:0] sltu_result;
wire [31:0] and_result;
wire [31:0] nor_result;
wire [31:0] or_result;
wire [31:0] xor_result;
wire [31:0] lui_result;
wire [31:0] sll_result; 
wire [63:0] sr64_result; 
wire [31:0] sr_result; 
wire [63:0] unsigned_prod_result;
wire [63:0] signed_prod_result;

// 32-bit adder
wire [31:0] adder_a;
wire [31:0] adder_b;
wire        adder_cin;
wire [31:0] adder_result;
wire        adder_cout;

assign adder_a   = alu_src1;
assign adder_b   = (op_sub | op_slt | op_sltu) ? ~alu_src2 : alu_src2;
assign adder_cin = (op_sub | op_slt | op_sltu) ? 1'b1      : 1'b0;
assign {adder_cout, adder_result} = adder_a + adder_b + adder_cin;

// ADD, SUB result
assign add_sub_result = adder_result;

// SLT result
assign slt_result[31:1] = 31'b0;
assign slt_result[0]    = (alu_src1[31] & ~alu_src2[31])
                        | ((alu_src1[31] ~^ alu_src2[31]) & adder_result[31]);

// SLTU result
assign sltu_result[31:1] = 31'b0;
assign sltu_result[0]    = ~adder_cout;

// bitwise operation
assign and_result = alu_src1 & alu_src2;
assign or_result  = alu_src1 | alu_src2;
assign nor_result = ~or_result;
assign xor_result = alu_src1 ^ alu_src2;
assign lui_result = {alu_src2[15:0], 16'b0};

// SLL result 
assign sll_result = alu_src2 << alu_src1[4:0];

// SRL, SRA result
assign sr64_result = {{32{op_sra & alu_src2[31]}}, alu_src2[31:0]} >> alu_src1[4:0];

assign sr_result   = sr64_result[31:0];

//MULT,MULTU result
assign unsigned_prod_result = alu_src1 * alu_src2;

assign signed_prod_result = $signed (alu_src1) * $signed (alu_src2);

// final result mux

assign alu_result   = ({32{op_add|op_sub}} & add_sub_result)
                     | ({32{op_slt       }} & slt_result)
                     | ({32{op_sltu      }} & sltu_result)
                     | ({32{op_and       }} & and_result)
                     | ({32{op_nor       }} & nor_result)
                     | ({32{op_or        }} & or_result)
                     | ({32{op_xor       }} & xor_result)
                     | ({32{op_lui       }} & lui_result)
                     | ({32{op_sll       }} & sll_result)
                     | ({32{op_srl|op_sra}} & sr_result)
                     | ({32{op_mul       }} & signed_prod_result[63:32])
                     | ({32{op_mul_n     }} & unsigned_prod_result[63:32])
                     | ({32{result_valid }} & result_data[63:32])
                     | ({32{result_valid_n }} & result_data_n[63:32]);


assign alu_result2  = ({32{op_mul       }} & signed_prod_result[31:0])
                    | ({32{op_mul_n     }} & unsigned_prod_result[31:0])
                    | ({32{result_valid }} & result_data[31:0])
                    | ({32{result_valid_n }} & result_data_n[31:0]);
endmodule
